/*****************************************************************************************
** 
**                               		北京交通大学                                     
**
**----------------------------------------------------------------------------------------
** 	文件名：			busComparator.v
** 	创建时间：		2015-8-18 10:00
** 	创建人员： 		赵秉贤
** 	文件描述：  		总线比较器源文件
** 
**----------------------------------------------------------------------------------------
** 	最后修改时间：	2015-8-18 10:00 
** 	最后修改人员：	赵秉贤
** 	版本号：	   	V1.0
** 	版本描述：		比较器基本逻辑梳理
**
*****************************************************************************************/

`timescale 1ps / 1ps

/*****************************************************************************************
**	模块名称:	busComparator()
**	模块功能:	比较器顶层模块
**	输入参数:	clk, rst
**	输出参数:	无
**	返回参数:	无
**	修改时间:	2015-8-18 10:12
*****************************************************************************************/
module busComparator(clk, rst);

input clk;
input rst;

always @(posedge clk or negedge clk) begin
	if(rst) begin
	
	end
	
	else begin
		/*初始化FIFO及输出状态*/
	end
end

endmodule



 